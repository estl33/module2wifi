-- nios_system.vhd

-- Generated using ACDS version 15.0 153

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system is
	port (
		bass_out_export     : out   std_logic_vector(3 downto 0);                     --     bass_out.export
		clk_clk             : in    std_logic                     := '0';             --          clk.clk
		hex0_1_export       : out   std_logic_vector(7 downto 0);                     --       hex0_1.export
		hex2_3_export       : out   std_logic_vector(7 downto 0);                     --       hex2_3.export
		hex4_5_export       : out   std_logic_vector(7 downto 0);                     --       hex4_5.export
		io_acknowledge      : in    std_logic                     := '0';             --           io.acknowledge
		io_irq              : in    std_logic                     := '0';             --             .irq
		io_address          : out   std_logic_vector(15 downto 0);                    --             .address
		io_bus_enable       : out   std_logic;                                        --             .bus_enable
		io_byte_enable      : out   std_logic_vector(1 downto 0);                     --             .byte_enable
		io_rw               : out   std_logic;                                        --             .rw
		io_write_data       : out   std_logic_vector(15 downto 0);                    --             .write_data
		io_read_data        : in    std_logic_vector(15 downto 0) := (others => '0'); --             .read_data
		lcd_data_DATA       : inout std_logic_vector(7 downto 0)  := (others => '0'); --     lcd_data.DATA
		lcd_data_ON         : out   std_logic;                                        --             .ON
		lcd_data_BLON       : out   std_logic;                                        --             .BLON
		lcd_data_EN         : out   std_logic;                                        --             .EN
		lcd_data_RS         : out   std_logic;                                        --             .RS
		lcd_data_RW         : out   std_logic;                                        --             .RW
		leds_export         : out   std_logic_vector(9 downto 0);                     --         leds.export
		push_buttons_export : in    std_logic_vector(2 downto 0)  := (others => '0'); -- push_buttons.export
		reset_reset_n       : in    std_logic                     := '0';             --        reset.reset_n
		sdram_addr          : out   std_logic_vector(12 downto 0);                    --        sdram.addr
		sdram_ba            : out   std_logic_vector(1 downto 0);                     --             .ba
		sdram_cas_n         : out   std_logic;                                        --             .cas_n
		sdram_cke           : out   std_logic;                                        --             .cke
		sdram_cs_n          : out   std_logic;                                        --             .cs_n
		sdram_dq            : inout std_logic_vector(15 downto 0) := (others => '0'); --             .dq
		sdram_dqm           : out   std_logic_vector(1 downto 0);                     --             .dqm
		sdram_ras_n         : out   std_logic;                                        --             .ras_n
		sdram_we_n          : out   std_logic;                                        --             .we_n
		sdram_clk_clk       : out   std_logic;                                        --    sdram_clk.clk
		sound_in_export     : in    std_logic_vector(15 downto 0) := (others => '0'); --     sound_in.export
		sound_out_export    : out   std_logic_vector(15 downto 0);                    --    sound_out.export
		switches_export     : in    std_logic_vector(9 downto 0)  := (others => '0'); --     switches.export
		treble_out_export   : out   std_logic_vector(3 downto 0);                     --   treble_out.export
		volume_out_export   : out   std_logic_vector(15 downto 0)                     --   volume_out.export
	);
end entity nios_system;

architecture rtl of nios_system is
	component nios_system_HEX0_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios_system_HEX0_1;

	component nios_system_PushButtons is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component nios_system_PushButtons;

	component nios_system_bass_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component nios_system_bass_out;

	component nios_system_character_lcd_0 is
		port (
			clk         : in    std_logic                    := 'X';             -- clk
			reset       : in    std_logic                    := 'X';             -- reset
			address     : in    std_logic                    := 'X';             -- address
			chipselect  : in    std_logic                    := 'X';             -- chipselect
			read        : in    std_logic                    := 'X';             -- read
			write       : in    std_logic                    := 'X';             -- write
			writedata   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                       -- waitrequest
			LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_ON      : out   std_logic;                                       -- export
			LCD_BLON    : out   std_logic;                                       -- export
			LCD_EN      : out   std_logic;                                       -- export
			LCD_RS      : out   std_logic;                                       -- export
			LCD_RW      : out   std_logic                                        -- export
		);
	end component nios_system_character_lcd_0;

	component nios_system_clocks is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component nios_system_clocks;

	component nios_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_system_jtag_uart_0;

	component nios_system_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component nios_system_leds;

	component nios_system_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(27 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic;                                        -- readra
			reset_req                             : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios_system_nios2_qsys_0;

	component nios_system_pot is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component nios_system_pot;

	component nios_system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_system_sdram;

	component nios_system_sound_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component nios_system_sound_in;

	component nios_system_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component nios_system_switches;

	component nios_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_system_timer_0;

	component nios_system_to_external_bus_bridge_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			avalon_address     : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			avalon_byteenable  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			avalon_chipselect  : in  std_logic                     := 'X';             -- chipselect
			avalon_read        : in  std_logic                     := 'X';             -- read
			avalon_write       : in  std_logic                     := 'X';             -- write
			avalon_writedata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avalon_readdata    : out std_logic_vector(15 downto 0);                    -- readdata
			avalon_waitrequest : out std_logic;                                        -- waitrequest
			avalon_irq         : out std_logic;                                        -- irq
			acknowledge        : in  std_logic                     := 'X';             -- export
			irq                : in  std_logic                     := 'X';             -- export
			address            : out std_logic_vector(15 downto 0);                    -- export
			bus_enable         : out std_logic;                                        -- export
			byte_enable        : out std_logic_vector(1 downto 0);                     -- export
			rw                 : out std_logic;                                        -- export
			write_data         : out std_logic_vector(15 downto 0);                    -- export
			read_data          : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component nios_system_to_external_bus_bridge_0;

	component nios_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                     : in  std_logic                     := 'X';             -- clk
			clocks_sys_clk_clk                                : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			sound_in_reset_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_data_master_address                  : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest              : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                     : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                    : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess              : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address           : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest       : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read              : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_instruction_master_readdatavalid     : out std_logic;                                        -- readdatavalid
			bass_out_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			bass_out_s1_write                                 : out std_logic;                                        -- write
			bass_out_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			bass_out_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			bass_out_s1_chipselect                            : out std_logic;                                        -- chipselect
			character_lcd_0_avalon_lcd_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			character_lcd_0_avalon_lcd_slave_write            : out std_logic;                                        -- write
			character_lcd_0_avalon_lcd_slave_read             : out std_logic;                                        -- read
			character_lcd_0_avalon_lcd_slave_readdata         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			character_lcd_0_avalon_lcd_slave_writedata        : out std_logic_vector(7 downto 0);                     -- writedata
			character_lcd_0_avalon_lcd_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			character_lcd_0_avalon_lcd_slave_chipselect       : out std_logic;                                        -- chipselect
			HEX0_1_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			HEX0_1_s1_write                                   : out std_logic;                                        -- write
			HEX0_1_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX0_1_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			HEX0_1_s1_chipselect                              : out std_logic;                                        -- chipselect
			HEX2_3_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			HEX2_3_s1_write                                   : out std_logic;                                        -- write
			HEX2_3_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX2_3_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			HEX2_3_s1_chipselect                              : out std_logic;                                        -- chipselect
			HEX4_5_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			HEX4_5_s1_write                                   : out std_logic;                                        -- write
			HEX4_5_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX4_5_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			HEX4_5_s1_chipselect                              : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write               : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			leds_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                     : out std_logic;                                        -- write
			leds_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                : out std_logic;                                        -- chipselect
			nios2_qsys_0_jtag_debug_module_address            : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_jtag_debug_module_write              : out std_logic;                                        -- write
			nios2_qsys_0_jtag_debug_module_read               : out std_logic;                                        -- read
			nios2_qsys_0_jtag_debug_module_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_jtag_debug_module_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess        : out std_logic;                                        -- debugaccess
			pot_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			pot_s1_write                                      : out std_logic;                                        -- write
			pot_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pot_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			pot_s1_chipselect                                 : out std_logic;                                        -- chipselect
			PushButtons_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			PushButtons_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_s1_address                                  : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                    : out std_logic;                                        -- write
			sdram_s1_read                                     : out std_logic;                                        -- read
			sdram_s1_readdata                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                               : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                            : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                              : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                               : out std_logic;                                        -- chipselect
			sound_in_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			sound_in_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sound_out_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			sound_out_s1_write                                : out std_logic;                                        -- write
			sound_out_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sound_out_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			sound_out_s1_chipselect                           : out std_logic;                                        -- chipselect
			switches_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                  : out std_logic;                                        -- write
			timer_0_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                             : out std_logic;                                        -- chipselect
			timer_1_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                                  : out std_logic;                                        -- write
			timer_1_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                             : out std_logic;                                        -- chipselect
			to_external_bus_bridge_0_avalon_slave_address     : out std_logic_vector(14 downto 0);                    -- address
			to_external_bus_bridge_0_avalon_slave_write       : out std_logic;                                        -- write
			to_external_bus_bridge_0_avalon_slave_read        : out std_logic;                                        -- read
			to_external_bus_bridge_0_avalon_slave_readdata    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			to_external_bus_bridge_0_avalon_slave_writedata   : out std_logic_vector(15 downto 0);                    -- writedata
			to_external_bus_bridge_0_avalon_slave_byteenable  : out std_logic_vector(1 downto 0);                     -- byteenable
			to_external_bus_bridge_0_avalon_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			to_external_bus_bridge_0_avalon_slave_chipselect  : out std_logic;                                        -- chipselect
			treble_out_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			treble_out_s1_write                               : out std_logic;                                        -- write
			treble_out_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			treble_out_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			treble_out_s1_chipselect                          : out std_logic                                         -- chipselect
		);
	end component nios_system_mm_interconnect_0;

	component nios_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component nios_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller;

	component nios_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_system_rst_controller_001;

	signal clocks_sys_clk_clk                                                  : std_logic;                     -- clocks:sys_clk_clk -> [HEX0_1:clk, HEX2_3:clk, HEX4_5:clk, PushButtons:clk, bass_out:clk, character_lcd_0:clk, irq_mapper:clk, irq_synchronizer:sender_clk, leds:clk, mm_interconnect_0:clocks_sys_clk_clk, nios2_qsys_0:clk, pot:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sound_in:clk, sound_out:clk, timer_0:clk, timer_1:clk, to_external_bus_bridge_0:clk, treble_out:clk]
	signal nios2_qsys_0_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_debugaccess                                : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_address                                    : std_logic_vector(27 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal nios2_qsys_0_data_master_read                                       : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_write                                      : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_writedata                                  : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal nios2_qsys_0_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                             : std_logic_vector(27 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                                : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal nios2_qsys_0_instruction_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect          : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata            : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest         : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write               : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect       : std_logic;                     -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_chipselect -> character_lcd_0:chipselect
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata         : std_logic_vector(7 downto 0);  -- character_lcd_0:readdata -> mm_interconnect_0:character_lcd_0_avalon_lcd_slave_readdata
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest      : std_logic;                     -- character_lcd_0:waitrequest -> mm_interconnect_0:character_lcd_0_avalon_lcd_slave_waitrequest
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_address -> character_lcd_0:address
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read             : std_logic;                     -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_read -> character_lcd_0:read
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write            : std_logic;                     -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_write -> character_lcd_0:write
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata        : std_logic_vector(7 downto 0);  -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_writedata -> character_lcd_0:writedata
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_chipselect  : std_logic;                     -- mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_chipselect -> to_external_bus_bridge_0:avalon_chipselect
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_readdata    : std_logic_vector(15 downto 0); -- to_external_bus_bridge_0:avalon_readdata -> mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_readdata
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_waitrequest : std_logic;                     -- to_external_bus_bridge_0:avalon_waitrequest -> mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_waitrequest
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_address     : std_logic_vector(14 downto 0); -- mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_address -> to_external_bus_bridge_0:avalon_address
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_read        : std_logic;                     -- mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_read -> to_external_bus_bridge_0:avalon_read
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_byteenable  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_byteenable -> to_external_bus_bridge_0:avalon_byteenable
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_write       : std_logic;                     -- mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_write -> to_external_bus_bridge_0:avalon_write
	signal mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_writedata   : std_logic_vector(15 downto 0); -- mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_writedata -> to_external_bus_bridge_0:avalon_writedata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata           : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest        : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess        : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read               : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write              : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal mm_interconnect_0_switches_s1_readdata                              : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_leds_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                                  : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                                     : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                 : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                              : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                  : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                     : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                            : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                    : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_hex0_1_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:HEX0_1_s1_chipselect -> HEX0_1:chipselect
	signal mm_interconnect_0_hex0_1_s1_readdata                                : std_logic_vector(31 downto 0); -- HEX0_1:readdata -> mm_interconnect_0:HEX0_1_s1_readdata
	signal mm_interconnect_0_hex0_1_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX0_1_s1_address -> HEX0_1:address
	signal mm_interconnect_0_hex0_1_s1_write                                   : std_logic;                     -- mm_interconnect_0:HEX0_1_s1_write -> mm_interconnect_0_hex0_1_s1_write:in
	signal mm_interconnect_0_hex0_1_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX0_1_s1_writedata -> HEX0_1:writedata
	signal mm_interconnect_0_hex4_5_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:HEX4_5_s1_chipselect -> HEX4_5:chipselect
	signal mm_interconnect_0_hex4_5_s1_readdata                                : std_logic_vector(31 downto 0); -- HEX4_5:readdata -> mm_interconnect_0:HEX4_5_s1_readdata
	signal mm_interconnect_0_hex4_5_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX4_5_s1_address -> HEX4_5:address
	signal mm_interconnect_0_hex4_5_s1_write                                   : std_logic;                     -- mm_interconnect_0:HEX4_5_s1_write -> mm_interconnect_0_hex4_5_s1_write:in
	signal mm_interconnect_0_hex4_5_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX4_5_s1_writedata -> HEX4_5:writedata
	signal mm_interconnect_0_hex2_3_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:HEX2_3_s1_chipselect -> HEX2_3:chipselect
	signal mm_interconnect_0_hex2_3_s1_readdata                                : std_logic_vector(31 downto 0); -- HEX2_3:readdata -> mm_interconnect_0:HEX2_3_s1_readdata
	signal mm_interconnect_0_hex2_3_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX2_3_s1_address -> HEX2_3:address
	signal mm_interconnect_0_hex2_3_s1_write                                   : std_logic;                     -- mm_interconnect_0:HEX2_3_s1_write -> mm_interconnect_0_hex2_3_s1_write:in
	signal mm_interconnect_0_hex2_3_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX2_3_s1_writedata -> HEX2_3:writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                               : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                                  : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                               : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                  : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_pushbuttons_s1_readdata                           : std_logic_vector(31 downto 0); -- PushButtons:readdata -> mm_interconnect_0:PushButtons_s1_readdata
	signal mm_interconnect_0_pushbuttons_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PushButtons_s1_address -> PushButtons:address
	signal mm_interconnect_0_sound_in_s1_readdata                              : std_logic_vector(31 downto 0); -- sound_in:readdata -> mm_interconnect_0:sound_in_s1_readdata
	signal mm_interconnect_0_sound_in_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sound_in_s1_address -> sound_in:address
	signal mm_interconnect_0_sound_out_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:sound_out_s1_chipselect -> sound_out:chipselect
	signal mm_interconnect_0_sound_out_s1_readdata                             : std_logic_vector(31 downto 0); -- sound_out:readdata -> mm_interconnect_0:sound_out_s1_readdata
	signal mm_interconnect_0_sound_out_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sound_out_s1_address -> sound_out:address
	signal mm_interconnect_0_sound_out_s1_write                                : std_logic;                     -- mm_interconnect_0:sound_out_s1_write -> mm_interconnect_0_sound_out_s1_write:in
	signal mm_interconnect_0_sound_out_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:sound_out_s1_writedata -> sound_out:writedata
	signal mm_interconnect_0_pot_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:pot_s1_chipselect -> pot:chipselect
	signal mm_interconnect_0_pot_s1_readdata                                   : std_logic_vector(31 downto 0); -- pot:readdata -> mm_interconnect_0:pot_s1_readdata
	signal mm_interconnect_0_pot_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pot_s1_address -> pot:address
	signal mm_interconnect_0_pot_s1_write                                      : std_logic;                     -- mm_interconnect_0:pot_s1_write -> mm_interconnect_0_pot_s1_write:in
	signal mm_interconnect_0_pot_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pot_s1_writedata -> pot:writedata
	signal mm_interconnect_0_treble_out_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:treble_out_s1_chipselect -> treble_out:chipselect
	signal mm_interconnect_0_treble_out_s1_readdata                            : std_logic_vector(31 downto 0); -- treble_out:readdata -> mm_interconnect_0:treble_out_s1_readdata
	signal mm_interconnect_0_treble_out_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:treble_out_s1_address -> treble_out:address
	signal mm_interconnect_0_treble_out_s1_write                               : std_logic;                     -- mm_interconnect_0:treble_out_s1_write -> mm_interconnect_0_treble_out_s1_write:in
	signal mm_interconnect_0_treble_out_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:treble_out_s1_writedata -> treble_out:writedata
	signal mm_interconnect_0_bass_out_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:bass_out_s1_chipselect -> bass_out:chipselect
	signal mm_interconnect_0_bass_out_s1_readdata                              : std_logic_vector(31 downto 0); -- bass_out:readdata -> mm_interconnect_0:bass_out_s1_readdata
	signal mm_interconnect_0_bass_out_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:bass_out_s1_address -> bass_out:address
	signal mm_interconnect_0_bass_out_s1_write                                 : std_logic;                     -- mm_interconnect_0:bass_out_s1_write -> mm_interconnect_0_bass_out_s1_write:in
	signal mm_interconnect_0_bass_out_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:bass_out_s1_writedata -> bass_out:writedata
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- to_external_bus_bridge_0:avalon_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver2_irq                                            : std_logic;                     -- timer_0:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                            : std_logic;                     -- timer_1:irq -> irq_mapper:receiver3_irq
	signal nios2_qsys_0_d_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_receiver_irq                                       : std_logic_vector(0 downto 0);  -- jtag_uart_0:av_irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [character_lcd_0:reset, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, to_external_bus_bridge_0:reset]
	signal nios2_qsys_0_jtag_debug_module_reset_reset                          : std_logic;                     -- nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:sound_in_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                                  : std_logic;                     -- rst_controller_002:reset_out -> clocks:ref_reset_reset
	signal rst_controller_003_reset_out_reset                                  : std_logic;                     -- rst_controller_003:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                           : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_hex0_1_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_hex0_1_s1_write:inv -> HEX0_1:write_n
	signal mm_interconnect_0_hex4_5_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_hex4_5_s1_write:inv -> HEX4_5:write_n
	signal mm_interconnect_0_hex2_3_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_hex2_3_s1_write:inv -> HEX2_3:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_sound_out_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_sound_out_s1_write:inv -> sound_out:write_n
	signal mm_interconnect_0_pot_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_pot_s1_write:inv -> pot:write_n
	signal mm_interconnect_0_treble_out_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_treble_out_s1_write:inv -> treble_out:write_n
	signal mm_interconnect_0_bass_out_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_bass_out_s1_write:inv -> bass_out:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [HEX0_1:reset_n, HEX2_3:reset_n, HEX4_5:reset_n, PushButtons:reset_n, leds:reset_n, nios2_qsys_0:reset_n, sdram:reset_n, timer_0:reset_n, timer_1:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [bass_out:reset_n, pot:reset_n, sound_in:reset_n, sound_out:reset_n, treble_out:reset_n]
	signal rst_controller_003_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> [jtag_uart_0:rst_n, switches:reset_n]

begin

	hex0_1 : component nios_system_HEX0_1
		port map (
			clk        => clocks_sys_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_hex0_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex0_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex0_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex0_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex0_1_s1_readdata,        --                    .readdata
			out_port   => hex0_1_export                                -- external_connection.export
		);

	hex2_3 : component nios_system_HEX0_1
		port map (
			clk        => clocks_sys_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_hex2_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex2_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex2_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex2_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex2_3_s1_readdata,        --                    .readdata
			out_port   => hex2_3_export                                -- external_connection.export
		);

	hex4_5 : component nios_system_HEX0_1
		port map (
			clk        => clocks_sys_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_hex4_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex4_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex4_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex4_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex4_5_s1_readdata,        --                    .readdata
			out_port   => hex4_5_export                                -- external_connection.export
		);

	pushbuttons : component nios_system_PushButtons
		port map (
			clk      => clocks_sys_clk_clk,                        --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_pushbuttons_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pushbuttons_s1_readdata, --                    .readdata
			in_port  => push_buttons_export                        -- external_connection.export
		);

	bass_out : component nios_system_bass_out
		port map (
			clk        => clocks_sys_clk_clk,                            --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_bass_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_bass_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_bass_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_bass_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_bass_out_s1_readdata,        --                    .readdata
			out_port   => bass_out_export                                -- external_connection.export
		);

	character_lcd_0 : component nios_system_character_lcd_0
		port map (
			clk         => clocks_sys_clk_clk,                                             --                clk.clk
			reset       => rst_controller_reset_out_reset,                                 --              reset.reset
			address     => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address(0),  --   avalon_lcd_slave.address
			chipselect  => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect,  --                   .chipselect
			read        => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read,        --                   .read
			write       => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write,       --                   .write
			writedata   => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest, --                   .waitrequest
			LCD_DATA    => lcd_data_DATA,                                                  -- external_interface.export
			LCD_ON      => lcd_data_ON,                                                    --                   .export
			LCD_BLON    => lcd_data_BLON,                                                  --                   .export
			LCD_EN      => lcd_data_EN,                                                    --                   .export
			LCD_RS      => lcd_data_RS,                                                    --                   .export
			LCD_RW      => lcd_data_RW                                                     --                   .export
		);

	clocks : component nios_system_clocks
		port map (
			ref_clk_clk        => clk_clk,                            --      ref_clk.clk
			ref_reset_reset    => rst_controller_002_reset_out_reset, --    ref_reset.reset
			sys_clk_clk        => clocks_sys_clk_clk,                 --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                      --    sdram_clk.clk
			reset_source_reset => open                                -- reset_source.reset
		);

	jtag_uart_0 : component nios_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_003_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_receiver_irq(0)                                 --               irq.irq
		);

	leds : component nios_system_leds
		port map (
			clk        => clocks_sys_clk_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_export                                -- external_connection.export
		);

	nios2_qsys_0 : component nios_system_nios2_qsys_0
		port map (
			clk                                   => clocks_sys_clk_clk,                                           --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                     --                   reset_n.reset_n
			d_address                             => nios2_qsys_0_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => nios2_qsys_0_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open,                                                         -- custom_instruction_master.readra
			reset_req                             => '0'                                                           --               (terminated)
		);

	pot : component nios_system_pot
		port map (
			clk        => clocks_sys_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_pot_s1_address,             --                  s1.address
			write_n    => mm_interconnect_0_pot_s1_write_ports_inv,     --                    .write_n
			writedata  => mm_interconnect_0_pot_s1_writedata,           --                    .writedata
			chipselect => mm_interconnect_0_pot_s1_chipselect,          --                    .chipselect
			readdata   => mm_interconnect_0_pot_s1_readdata,            --                    .readdata
			out_port   => volume_out_export                             -- external_connection.export
		);

	sdram : component nios_system_sdram
		port map (
			clk            => clocks_sys_clk_clk,                              --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sound_in : component nios_system_sound_in
		port map (
			clk      => clocks_sys_clk_clk,                           --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_sound_in_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_sound_in_s1_readdata,       --                    .readdata
			in_port  => sound_in_export                               -- external_connection.export
		);

	sound_out : component nios_system_pot
		port map (
			clk        => clocks_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_sound_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sound_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sound_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sound_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sound_out_s1_readdata,        --                    .readdata
			out_port   => sound_out_export                                -- external_connection.export
		);

	switches : component nios_system_switches
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,       --                    .readdata
			in_port  => switches_export                               -- external_connection.export
		);

	timer_0 : component nios_system_timer_0
		port map (
			clk        => clocks_sys_clk_clk,                           --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                      --   irq.irq
		);

	timer_1 : component nios_system_timer_0
		port map (
			clk        => clocks_sys_clk_clk,                           --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                      --   irq.irq
		);

	to_external_bus_bridge_0 : component nios_system_to_external_bus_bridge_0
		port map (
			clk                => clocks_sys_clk_clk,                                                  --                clk.clk
			reset              => rst_controller_reset_out_reset,                                      --              reset.reset
			avalon_address     => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_address,     --       avalon_slave.address
			avalon_byteenable  => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_byteenable,  --                   .byteenable
			avalon_chipselect  => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_chipselect,  --                   .chipselect
			avalon_read        => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_read,        --                   .read
			avalon_write       => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_write,       --                   .write
			avalon_writedata   => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_writedata,   --                   .writedata
			avalon_readdata    => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_readdata,    --                   .readdata
			avalon_waitrequest => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_waitrequest, --                   .waitrequest
			avalon_irq         => irq_mapper_receiver0_irq,                                            --          interrupt.irq
			acknowledge        => io_acknowledge,                                                      -- external_interface.export
			irq                => io_irq,                                                              --                   .export
			address            => io_address,                                                          --                   .export
			bus_enable         => io_bus_enable,                                                       --                   .export
			byte_enable        => io_byte_enable,                                                      --                   .export
			rw                 => io_rw,                                                               --                   .export
			write_data         => io_write_data,                                                       --                   .export
			read_data          => io_read_data                                                         --                   .export
		);

	treble_out : component nios_system_bass_out
		port map (
			clk        => clocks_sys_clk_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_treble_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_treble_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_treble_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_treble_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_treble_out_s1_readdata,        --                    .readdata
			out_port   => treble_out_export                                -- external_connection.export
		);

	mm_interconnect_0 : component nios_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                     => clk_clk,                                                             --                                  clk_0_clk.clk
			clocks_sys_clk_clk                                => clocks_sys_clk_clk,                                                  --                             clocks_sys_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset     => rst_controller_003_reset_out_reset,                                  --    jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                                      -- nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
			sound_in_reset_reset_bridge_in_reset_reset        => rst_controller_001_reset_out_reset,                                  --       sound_in_reset_reset_bridge_in_reset.reset
			nios2_qsys_0_data_master_address                  => nios2_qsys_0_data_master_address,                                    --                   nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest              => nios2_qsys_0_data_master_waitrequest,                                --                                           .waitrequest
			nios2_qsys_0_data_master_byteenable               => nios2_qsys_0_data_master_byteenable,                                 --                                           .byteenable
			nios2_qsys_0_data_master_read                     => nios2_qsys_0_data_master_read,                                       --                                           .read
			nios2_qsys_0_data_master_readdata                 => nios2_qsys_0_data_master_readdata,                                   --                                           .readdata
			nios2_qsys_0_data_master_write                    => nios2_qsys_0_data_master_write,                                      --                                           .write
			nios2_qsys_0_data_master_writedata                => nios2_qsys_0_data_master_writedata,                                  --                                           .writedata
			nios2_qsys_0_data_master_debugaccess              => nios2_qsys_0_data_master_debugaccess,                                --                                           .debugaccess
			nios2_qsys_0_instruction_master_address           => nios2_qsys_0_instruction_master_address,                             --            nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest       => nios2_qsys_0_instruction_master_waitrequest,                         --                                           .waitrequest
			nios2_qsys_0_instruction_master_read              => nios2_qsys_0_instruction_master_read,                                --                                           .read
			nios2_qsys_0_instruction_master_readdata          => nios2_qsys_0_instruction_master_readdata,                            --                                           .readdata
			nios2_qsys_0_instruction_master_readdatavalid     => nios2_qsys_0_instruction_master_readdatavalid,                       --                                           .readdatavalid
			bass_out_s1_address                               => mm_interconnect_0_bass_out_s1_address,                               --                                bass_out_s1.address
			bass_out_s1_write                                 => mm_interconnect_0_bass_out_s1_write,                                 --                                           .write
			bass_out_s1_readdata                              => mm_interconnect_0_bass_out_s1_readdata,                              --                                           .readdata
			bass_out_s1_writedata                             => mm_interconnect_0_bass_out_s1_writedata,                             --                                           .writedata
			bass_out_s1_chipselect                            => mm_interconnect_0_bass_out_s1_chipselect,                            --                                           .chipselect
			character_lcd_0_avalon_lcd_slave_address          => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address,          --           character_lcd_0_avalon_lcd_slave.address
			character_lcd_0_avalon_lcd_slave_write            => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write,            --                                           .write
			character_lcd_0_avalon_lcd_slave_read             => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read,             --                                           .read
			character_lcd_0_avalon_lcd_slave_readdata         => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata,         --                                           .readdata
			character_lcd_0_avalon_lcd_slave_writedata        => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata,        --                                           .writedata
			character_lcd_0_avalon_lcd_slave_waitrequest      => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest,      --                                           .waitrequest
			character_lcd_0_avalon_lcd_slave_chipselect       => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect,       --                                           .chipselect
			HEX0_1_s1_address                                 => mm_interconnect_0_hex0_1_s1_address,                                 --                                  HEX0_1_s1.address
			HEX0_1_s1_write                                   => mm_interconnect_0_hex0_1_s1_write,                                   --                                           .write
			HEX0_1_s1_readdata                                => mm_interconnect_0_hex0_1_s1_readdata,                                --                                           .readdata
			HEX0_1_s1_writedata                               => mm_interconnect_0_hex0_1_s1_writedata,                               --                                           .writedata
			HEX0_1_s1_chipselect                              => mm_interconnect_0_hex0_1_s1_chipselect,                              --                                           .chipselect
			HEX2_3_s1_address                                 => mm_interconnect_0_hex2_3_s1_address,                                 --                                  HEX2_3_s1.address
			HEX2_3_s1_write                                   => mm_interconnect_0_hex2_3_s1_write,                                   --                                           .write
			HEX2_3_s1_readdata                                => mm_interconnect_0_hex2_3_s1_readdata,                                --                                           .readdata
			HEX2_3_s1_writedata                               => mm_interconnect_0_hex2_3_s1_writedata,                               --                                           .writedata
			HEX2_3_s1_chipselect                              => mm_interconnect_0_hex2_3_s1_chipselect,                              --                                           .chipselect
			HEX4_5_s1_address                                 => mm_interconnect_0_hex4_5_s1_address,                                 --                                  HEX4_5_s1.address
			HEX4_5_s1_write                                   => mm_interconnect_0_hex4_5_s1_write,                                   --                                           .write
			HEX4_5_s1_readdata                                => mm_interconnect_0_hex4_5_s1_readdata,                                --                                           .readdata
			HEX4_5_s1_writedata                               => mm_interconnect_0_hex4_5_s1_writedata,                               --                                           .writedata
			HEX4_5_s1_chipselect                              => mm_interconnect_0_hex4_5_s1_chipselect,                              --                                           .chipselect
			jtag_uart_0_avalon_jtag_slave_address             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,             --              jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,               --                                           .write
			jtag_uart_0_avalon_jtag_slave_read                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                --                                           .read
			jtag_uart_0_avalon_jtag_slave_readdata            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,            --                                           .readdata
			jtag_uart_0_avalon_jtag_slave_writedata           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,           --                                           .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,         --                                           .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,          --                                           .chipselect
			leds_s1_address                                   => mm_interconnect_0_leds_s1_address,                                   --                                    leds_s1.address
			leds_s1_write                                     => mm_interconnect_0_leds_s1_write,                                     --                                           .write
			leds_s1_readdata                                  => mm_interconnect_0_leds_s1_readdata,                                  --                                           .readdata
			leds_s1_writedata                                 => mm_interconnect_0_leds_s1_writedata,                                 --                                           .writedata
			leds_s1_chipselect                                => mm_interconnect_0_leds_s1_chipselect,                                --                                           .chipselect
			nios2_qsys_0_jtag_debug_module_address            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,            --             nios2_qsys_0_jtag_debug_module.address
			nios2_qsys_0_jtag_debug_module_write              => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,              --                                           .write
			nios2_qsys_0_jtag_debug_module_read               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,               --                                           .read
			nios2_qsys_0_jtag_debug_module_readdata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,           --                                           .readdata
			nios2_qsys_0_jtag_debug_module_writedata          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,          --                                           .writedata
			nios2_qsys_0_jtag_debug_module_byteenable         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,         --                                           .byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest        => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest,        --                                           .waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess        => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess,        --                                           .debugaccess
			pot_s1_address                                    => mm_interconnect_0_pot_s1_address,                                    --                                     pot_s1.address
			pot_s1_write                                      => mm_interconnect_0_pot_s1_write,                                      --                                           .write
			pot_s1_readdata                                   => mm_interconnect_0_pot_s1_readdata,                                   --                                           .readdata
			pot_s1_writedata                                  => mm_interconnect_0_pot_s1_writedata,                                  --                                           .writedata
			pot_s1_chipselect                                 => mm_interconnect_0_pot_s1_chipselect,                                 --                                           .chipselect
			PushButtons_s1_address                            => mm_interconnect_0_pushbuttons_s1_address,                            --                             PushButtons_s1.address
			PushButtons_s1_readdata                           => mm_interconnect_0_pushbuttons_s1_readdata,                           --                                           .readdata
			sdram_s1_address                                  => mm_interconnect_0_sdram_s1_address,                                  --                                   sdram_s1.address
			sdram_s1_write                                    => mm_interconnect_0_sdram_s1_write,                                    --                                           .write
			sdram_s1_read                                     => mm_interconnect_0_sdram_s1_read,                                     --                                           .read
			sdram_s1_readdata                                 => mm_interconnect_0_sdram_s1_readdata,                                 --                                           .readdata
			sdram_s1_writedata                                => mm_interconnect_0_sdram_s1_writedata,                                --                                           .writedata
			sdram_s1_byteenable                               => mm_interconnect_0_sdram_s1_byteenable,                               --                                           .byteenable
			sdram_s1_readdatavalid                            => mm_interconnect_0_sdram_s1_readdatavalid,                            --                                           .readdatavalid
			sdram_s1_waitrequest                              => mm_interconnect_0_sdram_s1_waitrequest,                              --                                           .waitrequest
			sdram_s1_chipselect                               => mm_interconnect_0_sdram_s1_chipselect,                               --                                           .chipselect
			sound_in_s1_address                               => mm_interconnect_0_sound_in_s1_address,                               --                                sound_in_s1.address
			sound_in_s1_readdata                              => mm_interconnect_0_sound_in_s1_readdata,                              --                                           .readdata
			sound_out_s1_address                              => mm_interconnect_0_sound_out_s1_address,                              --                               sound_out_s1.address
			sound_out_s1_write                                => mm_interconnect_0_sound_out_s1_write,                                --                                           .write
			sound_out_s1_readdata                             => mm_interconnect_0_sound_out_s1_readdata,                             --                                           .readdata
			sound_out_s1_writedata                            => mm_interconnect_0_sound_out_s1_writedata,                            --                                           .writedata
			sound_out_s1_chipselect                           => mm_interconnect_0_sound_out_s1_chipselect,                           --                                           .chipselect
			switches_s1_address                               => mm_interconnect_0_switches_s1_address,                               --                                switches_s1.address
			switches_s1_readdata                              => mm_interconnect_0_switches_s1_readdata,                              --                                           .readdata
			timer_0_s1_address                                => mm_interconnect_0_timer_0_s1_address,                                --                                 timer_0_s1.address
			timer_0_s1_write                                  => mm_interconnect_0_timer_0_s1_write,                                  --                                           .write
			timer_0_s1_readdata                               => mm_interconnect_0_timer_0_s1_readdata,                               --                                           .readdata
			timer_0_s1_writedata                              => mm_interconnect_0_timer_0_s1_writedata,                              --                                           .writedata
			timer_0_s1_chipselect                             => mm_interconnect_0_timer_0_s1_chipselect,                             --                                           .chipselect
			timer_1_s1_address                                => mm_interconnect_0_timer_1_s1_address,                                --                                 timer_1_s1.address
			timer_1_s1_write                                  => mm_interconnect_0_timer_1_s1_write,                                  --                                           .write
			timer_1_s1_readdata                               => mm_interconnect_0_timer_1_s1_readdata,                               --                                           .readdata
			timer_1_s1_writedata                              => mm_interconnect_0_timer_1_s1_writedata,                              --                                           .writedata
			timer_1_s1_chipselect                             => mm_interconnect_0_timer_1_s1_chipselect,                             --                                           .chipselect
			to_external_bus_bridge_0_avalon_slave_address     => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_address,     --      to_external_bus_bridge_0_avalon_slave.address
			to_external_bus_bridge_0_avalon_slave_write       => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_write,       --                                           .write
			to_external_bus_bridge_0_avalon_slave_read        => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_read,        --                                           .read
			to_external_bus_bridge_0_avalon_slave_readdata    => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_readdata,    --                                           .readdata
			to_external_bus_bridge_0_avalon_slave_writedata   => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_writedata,   --                                           .writedata
			to_external_bus_bridge_0_avalon_slave_byteenable  => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_byteenable,  --                                           .byteenable
			to_external_bus_bridge_0_avalon_slave_waitrequest => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_waitrequest, --                                           .waitrequest
			to_external_bus_bridge_0_avalon_slave_chipselect  => mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_chipselect,  --                                           .chipselect
			treble_out_s1_address                             => mm_interconnect_0_treble_out_s1_address,                             --                              treble_out_s1.address
			treble_out_s1_write                               => mm_interconnect_0_treble_out_s1_write,                               --                                           .write
			treble_out_s1_readdata                            => mm_interconnect_0_treble_out_s1_readdata,                            --                                           .readdata
			treble_out_s1_writedata                           => mm_interconnect_0_treble_out_s1_writedata,                           --                                           .writedata
			treble_out_s1_chipselect                          => mm_interconnect_0_treble_out_s1_chipselect                           --                                           .chipselect
		);

	irq_mapper : component nios_system_irq_mapper
		port map (
			clk           => clocks_sys_clk_clk,             --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_qsys_0_d_irq_irq          --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => clocks_sys_clk_clk,                 --         sender_clk.clk
			receiver_reset => rst_controller_003_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	rst_controller : component nios_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clocks_sys_clk_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_001 : component nios_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clocks_sys_clk_clk,                 --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component nios_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => open,                                       --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_003 : component nios_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                                    --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_hex0_1_s1_write_ports_inv <= not mm_interconnect_0_hex0_1_s1_write;

	mm_interconnect_0_hex4_5_s1_write_ports_inv <= not mm_interconnect_0_hex4_5_s1_write;

	mm_interconnect_0_hex2_3_s1_write_ports_inv <= not mm_interconnect_0_hex2_3_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_sound_out_s1_write_ports_inv <= not mm_interconnect_0_sound_out_s1_write;

	mm_interconnect_0_pot_s1_write_ports_inv <= not mm_interconnect_0_pot_s1_write;

	mm_interconnect_0_treble_out_s1_write_ports_inv <= not mm_interconnect_0_treble_out_s1_write;

	mm_interconnect_0_bass_out_s1_write_ports_inv <= not mm_interconnect_0_bass_out_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of nios_system
